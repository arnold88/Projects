library verilog;
use verilog.vl_types.all;
entity md5testbench is
end md5testbench;
